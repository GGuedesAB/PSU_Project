** Profile: "SCHEMATIC1-simulation"  [ C:\Users\Gustavo\Dropbox\UFMG\6 Periodo\Lab ELT1\Projetos\rectificationstage-pspicefiles\schematic1\simulation.sim ] 

** Creating circuit file "simulation.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../rectificationstage-PSpiceFiles/RECTIFICATIONSTAGE.lib" 
* From [PSPICE NETLIST] section of C:\Users\Gustavo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 10u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
